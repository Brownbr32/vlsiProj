/home/bbrown/IC_CAD/CADENCE/PVS_LVS/netlist